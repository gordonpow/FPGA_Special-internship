library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FPGA_VGA is
    Port (
        i_clk       : in STD_LOGIC;
        i_rst       : in STD_LOGIC;
        i_led_state : in STD_LOGIC_VECTOR(7 downto 0);
        hsync       : out STD_LOGIC;
        vsync       : out STD_LOGIC;
        red         : out STD_LOGIC_VECTOR (3 downto 0);
        green       : out STD_LOGIC_VECTOR (3 downto 0);
        blue        : out STD_LOGIC_VECTOR (3 downto 0)
    );
end FPGA_VGA;

architecture Behavioral of FPGA_VGA is

    -- VGA 640x480 @ 60 Hz �Ѽ�
    constant hRez        : integer := 640;
    constant hStartSync  : integer := 656;
    constant hEndSync    : integer := 752;
    constant hMaxCount   : integer := 800;

    constant vRez        : integer := 480;
    constant vStartSync  : integer := 490;
    constant vEndSync    : integer := 492;
    constant vMaxCount   : integer := 525;

    signal hCount : integer := 0;
    signal vCount : integer := 0;
    signal div    : STD_LOGIC_VECTOR(60 downto 0);
    signal vga_clk: STD_LOGIC;
    
    -- ø�Ϭ����T��
    signal slot_index : integer range 0 to 7;
    signal slot_center_x : integer;
    signal diff_x : integer;
    signal diff_y : integer;
    
    -- ��Υb�|���� (R=25, R^2=625) �y�L�Y�p�@�I�קK�H�b�@�_
    constant ball_r_sq : integer := 625; 
    -- ��� Y �y��
    constant ball_center_y : integer := 240;

begin
    -- ���� VGA Clock
    process(i_clk, i_rst)
    begin
        if i_rst = '1' then 
            div <= (others => '0');
        elsif rising_edge(i_clk) then 
            div <= div + 1;
        end if;
    end process;
    vga_clk <= div(1);

    -- �����P�����p�ƾ�
    process(vga_clk)
    begin
        if rising_edge(vga_clk) then
            if hCount = hMaxCount - 1 then
                hCount <= 0;
                if vCount = vMaxCount - 1 then
                    vCount <= 0;
                else
                    vCount <= vCount + 1;
                end if;
            else
                hCount <= hCount + 1;
            end if;
        end if;
    end process;

    -- �P�B�T��
    hsync <= '0' when (hCount >= hStartSync and hCount < hEndSync) else '1';
    vsync <= '0' when (vCount >= vStartSync and vCount < vEndSync) else '1';

    -- [�֤��޿�ץ�]
    -- 1. �ѨM�h���O���G�G���p���@�y�y�СA�ӬO�p���e�����ݩ���@�� LED ���u���Ұϡv�C
    -- 2. �ѨM��V�ۤϡG�����վ� bit ���� (Slot 0 ���� Bit 0, Slot 7 ���� Bit 7)�C
    
    process(hCount, vCount, i_led_state)
        variable current_bit_active : boolean;
        variable dx : integer;
        variable dy : integer;
    begin        
        if (hCount < hRez and vCount < vRez) then
            
            -- �p��ثe���y�u�b���@�Ӱ϶� (0~7)
            -- �C�Ӱ϶��e 80 pixel
            if hCount < 640 then
                slot_index <= hCount / 80;
            else
                slot_index <= 0;
            end if;

            -- �p��Ӱ϶������� X �I
            -- Slot 0 ����=40, Slot 1 ����=120... ����: index*80 + 40
            slot_center_x <= (hCount / 80) * 80 + 40;

            -- ���o�۹�Z�� (������ȷ���)
            if hCount > slot_center_x then
                dx := hCount - slot_center_x;
            else
                dx := slot_center_x - hCount;
            end if;

            if vCount > ball_center_y then
                dy := vCount - ball_center_y;
            else
                dy := ball_center_y - vCount;
            end if;

            -- �P�_�ثe�϶������� LED �O�_�G�_
            -- �i�o�̭ץ��F��V�j�G
            -- Slot 0 (�ù��̥�) ���� i_led_state(0)
            -- Slot 7 (�ù��̥k) ���� i_led_state(7)
            -- �p�G�o�٬O�Ϫ��A�Ч令 i_led_state(7 - (hCount / 80))
            if (hCount < 640) then
                if i_led_state(hCount / 80) = '1' then
                    current_bit_active := true;
                else
                    current_bit_active := false;
                end if;
            else
                current_bit_active := false;
            end if;

            -- ø���޿�
            -- �p�G 1. �ثe�����b��νd�� �B 2. �Ӧ�m��LED�O�G��
            if (current_bit_active) and ((dx*dx + dy*dy) < ball_r_sq) then
                -- �G�O (����)
                red   <= "1111";
                green <= "1111";
                blue  <= "0000";
            else
                -- �I�� (�`��)
                red   <= "0000";
                green <= "0000";
                blue  <= "0010";
            end if;
            
        else
            -- Blanking
            red   <= "0000";
            green <= "0000";
            blue  <= "0000";
        end if;
    end process;

end Behavioral;